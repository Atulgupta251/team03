module top_module(input [63:0] a, input[47:0] key, output [63:0] b);
    wire [63:0] x,y;
    wire [47:0] z,w;
    wire [31:0] v,u;
    bitpermute IP(a,x);
    y[63:32] = x[31:0];
    expansion E(a[31:0], z);
    assign w = z ^ key;
    S1Box S1(w[47:42], v[31:28]);
    S2Box S2(w[41:36], v[27:24]);
    S3Box S3(w[35:30], v[23:20]);
    S4Box S4(w[29:24], v[19:16]);
    S5Box S5(w[23:18], v[15:12]);
    S6Box S6(w[17:12], v[11: 8]);
    S7Box S7(w[11: 6], v[ 7: 4]);
    S8Box S8(w[ 5: 0], v[ 3: 0]);
    
    permute(v,u);
    assign y[31:0] = x[63:31] ^ u ;
    
    inversebitpermute IP_Inverse(y,b);
    
endmodule
   
module S1Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
    b[0][0] = 4'b1110;
    b[0][1] = 4'b0100;
    b[0][2] = 4'b1101;
    b[0][3] = 4'b0001;
    b[0][4] = 4'b0010;
    b[0][5] = 4'b1111;
    b[0][6] = 4'b1011;
    b[0][7] = 4'b1000;
    b[0][8] = 4'b0011;
    b[0][9] = 4'b1010;
    b[0][10] = 4'b0110;
    b[0][11] = 4'b1100;
    b[0][12] = 4'b0101;
    b[0][13] = 4'b1001;
    b[0][14] = 4'b0000;
    b[0][15] = 4'b0111;
            
    b[1][0] = 4'b0000;
    b[1][1] = 4'b1111;
    b[1][2] = 4'b0111;
    b[1][3] = 4'b0100;
    b[1][4] = 4'b1110;
    b[1][5] = 4'b0010;
    b[1][6] = 4'b1101;
    b[1][7] = 4'b0001;
    b[1][8] = 4'b1010;
    b[1][9] = 4'b0110;
    b[1][10] = 4'b1100;
    b[1][11] = 4'b1011;
    b[1][12] = 4'b1001;
    b[1][13] = 4'b0101;
    b[1][14] = 4'b0011;
    b[1][15] = 4'b1000;
            
    b[2][0] = 4'b0100;
    b[2][1] = 4'b0001;
    b[2][2] = 4'b1110;
    b[2][3] = 4'b1000;
    b[2][4] = 4'b1101;
    b[2][5] = 4'b0110;
    b[2][6] = 4'b0010;
    b[2][7] = 4'b1011;
    b[2][8] = 4'b1111;
    b[2][9] = 4'b1100;
    b[2][10] = 4'b1001;
    b[2][11] = 4'b0111;
    b[2][12] = 4'b0011;
    b[2][13] = 4'b1100;
    b[2][14] = 4'b0101;
    b[2][15] = 4'b0000;
            
    b[3][0] = 4'b1111;
    b[3][1] = 4'b1100;
    b[3][2] = 4'b1000;
    b[3][3] = 4'b0010;
    b[3][4] = 4'b0100;
    b[3][5] = 4'b1001;
    b[3][6] = 4'b0001;
    b[3][7] = 4'b0111;
    b[3][8] = 4'b0101;
    b[3][9] = 4'b1101;
    b[3][10] = 4'b0011;
    b[3][11] = 4'b1110;
    b[3][12] = 4'b1100;
    b[3][13] = 4'b0000;
    b[3][14] = 4'b0110;
    b[3][15] = 4'b1101;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S2Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
        b[0][0] = 4'b1111;
        b[0][1] = 4'b0001;
        b[0][2] = 4'b1000;
        b[0][3] = 4'b1110;
        b[0][4] = 4'b0110;
        b[0][5] = 4'b1011;
        b[0][6] = 4'b0011;
        b[0][7] = 4'b0100;
        b[0][8] = 4'b1001
        b[0][9] = 4'b0111;
        b[0][10] = 4'b0010;
        b[0][11] = 4'b1101;
        b[0][12] = 4'b1101;
        b[0][13] = 4'b0000;
        b[0][14] = 4'b0101;
        b[0][15] = 4'b1010;
            
        b[1][0] = 4'b0011;
        b[1][1] = 4'b1101;
        b[1][2] = 4'b0100;
        b[1][3] = 4'b0111;
        b[1][4] = 4'b1111;
        b[1][5] = 4'b0010;
        b[1][6] = 4'b1000;
        b[1][7] = 4'b1110;
        b[1][8] = 4'b1100;
        b[1][9] = 4'b0000;
        b[1][10] = 4'b0001;
        b[1][11] = 4'b1100;
        b[1][12] = 4'b0110;
        b[1][13] = 4'b1001;
        b[1][14] = 4'b1101;
        b[1][15] = 4'b0101;
            
        b[2][0] = 4'b0000;
        b[2][1] = 4'b1110;
        b[2][2] = 4'b0111;
        b[2][3] = 4'b1101;
        b[2][4] = 4'b1100;
        b[2][5] = 4'b0100;
        b[2][6] = 4'b1101;
        b[2][7] = 4'b0001;
        b[2][8] = 4'b0101;
        b[2][9] = 4'b1000;
        b[2][10] = 4'b1100;
        b[2][11] = 4'b0110;
        b[2][12] = 4'b1001;
        b[2][13] = 4'b0011;
        b[2][14] = 4'b0010;
        b[2][15] = 4'b1111;
            
        b[3][0] = 4'b1101;
        b[3][1] = 4'b1000;
        b[3][2] = 4'b1100;
        b[3][3] = 4'b0001;
        b[3][4] = 4'b0011;
        b[3][5] = 4'b1111;
        b[3][6] = 4'b0100;
        b[3][7] = 4'b0010;
        b[3][8] = 4'b1101;
        b[3][9] = 4'b0110;
        b[3][10] = 4'b0111;
        b[3][11] = 4'b1100;
        b[3][12] = 4'b0000;
        b[3][13] = 4'b0101;
        b[3][14] = 4'b1110;
        b[3][15] = 4'b1001;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S3Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
        b[0][0] = 4'b1100;
        b[0][1] = 4'b0000;
        b[0][2] = 4'b1001;
        b[0][3] = 4'b1110;
        b[0][4] = 4'b0110;
        b[0][5] = 4'b0011;
        b[0][6] = 4'b1111;
        b[0][7] = 4'b0101;
        b[0][8] = 4'b0001
        b[0][9] = 4'b1101;
        b[0][10] = 4'b1100;
        b[0][11] = 4'b0111;
        b[0][12] = 4'b1011;
        b[0][13] = 4'b0100;
        b[0][14] = 4'b0010;
        b[0][15] = 4'b1000;
            
        b[1][0] = 4'b1101;
        b[1][1] = 4'b0111;
        b[1][2] = 4'b0000;
        b[1][3] = 4'b1001;
        b[1][4] = 4'b0011;
        b[1][5] = 4'b0100;
        b[1][6] = 4'b0110;
        b[1][7] = 4'b1100;
        b[1][8] = 4'b0010;
        b[1][9] = 4'b1000;
        b[1][10] = 4'b0101;
        b[1][11] = 4'b1110;
        b[1][12] = 4'b1100;
        b[1][13] = 4'b1011;
        b[1][14] = 4'b1111;
        b[1][15] = 4'b0001;
            
        b[2][0] = 4'b1101;
        b[2][1] = 4'b0110;
        b[2][2] = 4'b0100;
        b[2][3] = 4'b1001;
        b[2][4] = 4'b1000;
        b[2][5] = 4'b1111;
        b[2][6] = 4'b0011;
        b[2][7] = 4'b0000;
        b[2][8] = 4'b1011;
        b[2][9] = 4'b0001;
        b[2][10] = 4'b0010;
        b[2][11] = 4'b1100;
        b[2][12] = 4'b0101;
        b[2][13] = 4'b1100;
        b[2][14] = 4'b1110;
        b[2][15] = 4'b0111;
            
        b[3][0] = 4'b0001;
        b[3][1] = 4'b1100;
        b[3][2] = 4'b1101;
        b[3][3] = 4'b0000;
        b[3][4] = 4'b0110;
        b[3][5] = 4'b1001;
        b[3][6] = 4'b1000;
        b[3][7] = 4'b0111;
        b[3][8] = 4'b0100;
        b[3][9] = 4'b1111;
        b[3][10] = 4'b1110;
        b[3][11] = 4'b0011;
        b[3][12] = 4'b1011;
        b[3][13] = 4'b0101;
        b[3][14] = 4'b0010;
        b[3][15] = 4'b1100;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S4Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
        b[0][0] = 4'b0111;
        b[0][1] = 4'b1101;
        b[0][2] = 4'b1110;
        b[0][3] = 4'b0011;
        b[0][4] = 4'b0000;
        b[0][5] = 4'b0110;
        b[0][6] = 4'b1001;
        b[0][7] = 4'b1010;
        b[0][8] = 4'b0001
        b[0][9] = 4'b0010;
        b[0][10] = 4'b1000;
        b[0][11] = 4'b0101;
        b[0][12] = 4'b1011;
        b[0][13] = 4'b1100;
        b[0][14] = 4'b0100;
        b[0][15] = 4'b1111;
            
        b[1][0] = 4'b1101;
        b[1][1] = 4'b1000;
        b[1][2] = 4'b1011;
        b[1][3] = 4'b0101;
        b[1][4] = 4'b0110;
        b[1][5] = 4'b1111;
        b[1][6] = 4'b0000;
        b[1][7] = 4'b0011;
        b[1][8] = 4'b0100;
        b[1][9] = 4'b0111;
        b[1][10] = 4'b0010;
        b[1][11] = 4'b1100;
        b[1][12] = 4'b0001;
        b[1][13] = 4'b1010;
        b[1][14] = 4'b1110;
        b[1][15] = 4'b1001;
            
        b[2][0] = 4'b1010;
        b[2][1] = 4'b0110;
        b[2][2] = 4'b1001;
        b[2][3] = 4'b0000;
        b[2][4] = 4'b1100;
        b[2][5] = 4'b1011;
        b[2][6] = 4'b0111;
        b[2][7] = 4'b1101;
        b[2][8] = 4'b1111;
        b[2][9] = 4'b0001;
        b[2][10] = 4'b0011;
        b[2][11] = 4'b1110;
        b[2][12] = 4'b0101;
        b[2][13] = 4'b0010;
        b[2][14] = 4'b1000;
        b[2][15] = 4'b0100;
            
        b[3][0] = 4'b0011;
        b[3][1] = 4'b1111;
        b[3][2] = 4'b0000;
        b[3][3] = 4'b0110;
        b[3][4] = 4'b1010;
        b[3][5] = 4'b0001;
        b[3][6] = 4'b1101;
        b[3][7] = 4'b1000;
        b[3][8] = 4'b1001;
        b[3][9] = 4'b0100;
        b[3][10] = 4'b0101;
        b[3][11] = 4'b1011;
        b[3][12] = 4'b1100;
        b[3][13] = 4'b0111;
        b[3][14] = 4'b0010;
        b[3][15] = 4'b1110;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S5Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
    b[0][0] = 4'b0010;
    b[0][1] = 4'b1100;
    b[0][2] = 4'b0100;
    b[0][3] = 4'b0001;
    b[0][4] = 4'b0111;
    b[0][5] = 4'b1010;
    b[0][6] = 4'b1011;
    b[0][7] = 4'b0110;
    b[0][8] = 4'b1000;
    b[0][9] = 4'b0101;
    b[0][10] = 4'b0011;
    b[0][11] = 4'b1011;
    b[0][12] = 4'b1101;
    b[0][13] = 4'b0000;
    b[0][14] = 4'b1110;
    b[0][15] = 4'b1001;
            
    b[1][0] = 4'b1110;
    b[1][1] = 4'b1011;
    b[1][2] = 4'b0010;
    b[1][3] = 4'b1100;
    b[1][4] = 4'b0100;
    b[1][5] = 4'b0111;
    b[1][6] = 4'b1101;
    b[1][7] = 4'b0001;
    b[1][8] = 4'b0101;
    b[1][9] = 4'b0000;
    b[1][10] = 4'b1111;
    b[1][11] = 4'b1010;
    b[1][12] = 4'b0011;
    b[1][13] = 4'b1001;
    b[1][14] = 4'b1000;
    b[1][15] = 4'b0110;
            
    b[2][0] = 4'b0100;
    b[2][1] = 4'b0010;
    b[2][2] = 4'b0001;
    b[2][3] = 4'b1011;
    b[2][4] = 4'b1010;
    b[2][5] = 4'b1101;
    b[2][6] = 4'b0111;
    b[2][7] = 4'b1000;
    b[2][8] = 4'b1111;
    b[2][9] = 4'b1001;
    b[2][10] = 4'b1100;
    b[2][11] = 4'b0101;
    b[2][12] = 4'b0110;
    b[2][13] = 4'b0011;
    b[2][14] = 4'b0000;
    b[2][15] = 4'b1110;
            
    b[3][0] = 4'b1011;
    b[3][1] = 4'b1000;
    b[3][2] = 4'b1100;
    b[3][3] = 4'b0111;
    b[3][4] = 4'b0001;
    b[3][5] = 4'b1110;
    b[3][6] = 4'b0010;
    b[3][7] = 4'b1101;
    b[3][8] = 4'b0110;
    b[3][9] = 4'b1111;
    b[3][10] = 4'b0000;
    b[3][11] = 4'b1001;
    b[3][12] = 4'b1010;
    b[3][13] = 4'b0100;
    b[3][14] = 4'b0101;
    b[3][15] = 4'b0011;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S6Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
    b[0][0] = 4'b1100;
    b[0][1] = 4'b0001;
    b[0][2] = 4'b1010;
    b[0][3] = 4'b1111;
    b[0][4] = 4'b1001;
    b[0][5] = 4'b0010;
    b[0][6] = 4'b0110;
    b[0][7] = 4'b1000;
    b[0][8] = 4'b0000;
    b[0][9] = 4'b1101;
    b[0][10] = 4'b0011;
    b[0][11] = 4'b0100;
    b[0][12] = 4'b1110;
    b[0][13] = 4'b0111;
    b[0][14] = 4'b0101;
    b[0][15] = 4'b1011;
            
    b[1][0] = 4'b1010;
    b[1][1] = 4'b1111;
    b[1][2] = 4'b0100;
    b[1][3] = 4'b0010;
    b[1][4] = 4'b0111;
    b[1][5] = 4'b1100;
    b[1][6] = 4'b1001;
    b[1][7] = 4'b0101;
    b[1][8] = 4'b0110;
    b[1][9] = 4'b0001;
    b[1][10] = 4'b1101;
    b[1][11] = 4'b1110;
    b[1][12] = 4'b0000;
    b[1][13] = 4'b1011;
    b[1][14] = 4'b0011;
    b[1][15] = 4'b1011;
            
    b[2][0] = 4'b1001;
    b[2][1] = 4'b1110;
    b[2][2] = 4'b1111;
    b[2][3] = 4'b0101;
    b[2][4] = 4'b0010;
    b[2][5] = 4'b1000;
    b[2][6] = 4'b1100;
    b[2][7] = 4'b0011;
    b[2][8] = 4'b0111;
    b[2][9] = 4'b0000;
    b[2][10] = 4'b0100;
    b[2][11] = 4'b1010;
    b[2][12] = 4'b0001;
    b[2][13] = 4'b1101;
    b[2][14] = 4'b1011;
    b[2][15] = 4'b0110;
            
    b[3][0] = 4'b0100;
    b[3][1] = 4'b0011;
    b[3][2] = 4'b0010;
    b[3][3] = 4'b1100;
    b[3][4] = 4'b1001;
    b[3][5] = 4'b0101;
    b[3][6] = 4'b1111;
    b[3][7] = 4'b1010;
    b[3][8] = 4'b1011;
    b[3][9] = 4'b1110;
    b[3][10] = 4'b0001;
    b[3][11] = 4'b0111;
    b[3][12] = 4'b1010;
    b[3][13] = 4'b0000;
    b[3][14] = 4'b1000;
    b[3][15] = 4'b1101;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S7Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
    b[0][0] = 4'b0100;
    b[0][1] = 4'b1011;
    b[0][2] = 4'b0010;
    b[0][3] = 4'b1110;
    b[0][4] = 4'b1111;
    b[0][5] = 4'b0000;
    b[0][6] = 4'b1000;
    b[0][7] = 4'b1101;
    b[0][8] = 4'b0011;
    b[0][9] = 4'b1100;
    b[0][10] = 4'b1001;
    b[0][11] = 4'b0111;
    b[0][12] = 4'b0101;
    b[0][13] = 4'b1010;
    b[0][14] = 4'b0110;
    b[0][15] = 4'b0001;
            
    b[1][0] = 4'b1101;
    b[1][1] = 4'b0000;
    b[1][2] = 4'b1011;
    b[1][3] = 4'b0111;
    b[1][4] = 4'b0100;
    b[1][5] = 4'b1001;
    b[1][6] = 4'b0001;
    b[1][7] = 4'b1010;
    b[1][8] = 4'b1110;
    b[1][9] = 4'b0011;
    b[1][10] = 4'b0101;
    b[1][11] = 4'b1100;
    b[1][12] = 4'b0010;
    b[1][13] = 4'b1111;
    b[1][14] = 4'b1000;
    b[1][15] = 4'b0110;
            
    b[2][0] = 4'b0001;
    b[2][1] = 4'b0100;
    b[2][2] = 4'b1101;
    b[2][3] = 4'b1101;
    b[2][4] = 4'b1100;
    b[2][5] = 4'b0011;
    b[2][6] = 4'b0111;
    b[2][7] = 4'b1110;
    b[2][8] = 4'b1010;
    b[2][9] = 4'b1111;
    b[2][10] = 4'b0110;
    b[2][11] = 4'b1000;
    b[2][12] = 4'b0000;
    b[2][13] = 4'b0101;
    b[2][14] = 4'b1001;
    b[2][15] = 4'b0010;
            
    b[3][0] = 4'b0110;
    b[3][1] = 4'b1011;
    b[3][2] = 4'b1101;
    b[3][3] = 4'b1000;
    b[3][4] = 4'b0001;
    b[3][5] = 4'b0100;
    b[3][6] = 4'b1010;
    b[3][7] = 4'b0111;
    b[3][8] = 4'b1001;
    b[3][9] = 4'b0101;
    b[3][10] = 4'b0000;
    b[3][11] = 4'b1111;
    b[3][12] = 4'b1110;
    b[3][13] = 4'b0010;
    b[3][14] = 4'b0011;
    b[3][15] = 4'b1100;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule

module S8Box(input [5:0] a, output [3:0] out);
    reg [3:0] b[0:3][0:15];
    initial begin
    b[0][0] = 4'b1101;
    b[0][1] = 4'b0010;
    b[0][2] = 4'b1000;
    b[0][3] = 4'b0100;
    b[0][4] = 4'b0110;
    b[0][5] = 4'b1111;
    b[0][6] = 4'b1011;
    b[0][7] = 4'b0001;
    b[0][8] = 4'b1010;
    b[0][9] = 4'b1001;
    b[0][10] = 4'b0011;
    b[0][11] = 4'b1110;
    b[0][12] = 4'b0101;
    b[0][13] = 4'b0000;
    b[0][14] = 4'b1100;
    b[0][15] = 4'b0111;
            
    b[1][0] = 4'b0001;
    b[1][1] = 4'b1111;
    b[1][2] = 4'b1101;
    b[1][3] = 4'b1000;
    b[1][4] = 4'b0100;
    b[1][5] = 4'b0011;
    b[1][6] = 4'b0111;
    b[1][7] = 4'b0100;
    b[1][8] = 4'b1100;
    b[1][9] = 4'b0101;
    b[1][10] = 4'b0110;
    b[1][11] = 4'b1011;
    b[1][12] = 4'b1010;
    b[1][13] = 4'b1110;
    b[1][14] = 4'b1001;
    b[1][15] = 4'b0010;
            
    b[2][0] = 4'b0111;
    b[2][1] = 4'b1011;
    b[2][2] = 4'b0100;
    b[2][3] = 4'b0001;
    b[2][4] = 4'b1001;
    b[2][5] = 4'b1100;
    b[2][6] = 4'b1110;
    b[2][7] = 4'b0010;
    b[2][8] = 4'b0000;
    b[2][9] = 4'b0110;
    b[2][10] = 4'b1010;
    b[2][11] = 4'b1010;
    b[2][12] = 4'b1111;
    b[2][13] = 4'b0011;
    b[2][14] = 4'b0101;
    b[2][15] = 4'b1000;
            
    b[3][0] = 4'b0010;
    b[3][1] = 4'b0001;
    b[3][2] = 4'b1110;
    b[3][3] = 4'b0111;
    b[3][4] = 4'b0100;
    b[3][5] = 4'b1010;
    b[3][6] = 4'b1000;
    b[3][7] = 4'b1101;
    b[3][8] = 4'b1111;
    b[3][9] = 4'b1100;
    b[3][10] = 4'b1001;
    b[3][11] = 4'b1001;
    b[3][12] = 4'b0011;
    b[3][13] = 4'b0101;
    b[3][14] = 4'b0110;
    b[3][15] = 4'b1011;
    end
    wire [3:0] col = a[4:1];
    wire [1:0] row = {a[5],a[0]};
    integer r,c;
    assign r = row;
    assign c = col;
    
    assign out = b[r][c];
    
endmodule




module Expansion(input [31:0] a, output [47:0] b);
    assign b ={a[31], a[ 0], a[ 1], a[ 2], a[ 3], a[ 4],
               a[ 3], a[ 4], a[ 5], a[ 6], a[ 7], a[ 8],
               a[ 7], a[ 8], a[ 9], a[10], a[11], a[12],
               a[11], a[16], a[13], a[14], a[15], a[16],
               a[15], a[20], a[17], a[18], a[19], a[20],
               a[19], a[24], a[21], a[22], a[23], a[24],
               a[23], a[28], a[25], a[26], a[27], a[28],
               a[27], a[32], a[29], a[30], a[31], a[ 0] };
endmodule





module bitpermute(input [63:0]a,output [63:0]b);
b[0]=a[5];b[1]=a[10];b[2]=a[15];b[3]=a[20];b[4]=a[25];b[5]=a[30];b[6]=a[35];b[7]=a[40];b[8]=a[45];b[9]=a[50];b[10]=a[55];b[11]=a[60];b[12]=a[1];b[13]=a[6];b[14]=a[11];b[15]=a[16];b[16]=a[21];b[17]=a[26];b[18]=a[31];b[19]=a[36];b[20]=a[41];b[21]=a[46];b[22]=a[51];b[23]=a[56];b[24]=a[61];b[25]=a[2];b[26]=a[7];b[27]=a[12];b[28]=a[17];b[29]=a[22];b[30]=a[27];b[31]=a[32];b[32]=a[37];b[33]=a[42];b[34]=a[47];b[35]=a[52];b[36]=a[57];b[37]=a[62];b[38]=a[3];b[39]=a[8];b[40]=a[13];b[41]=a[18];b[42]=a[23];b[43]=a[28];b[44]=a[33];b[45]=a[38];b[46]=a[43];b[47]=a[48];b[48]=a[53];b[49]=a[58];b[50]=a[63];b[51]=a[4];b[52]=a[9];b[53]=a[14];b[54]=a[19];b[55]=a[24];b[56]=a[29];b[57]=a[34];b[58]=a[39];b[59]=a[44];b[60]=a[49];b[61]=a[54];b[62]=a[59];b[63]=a[0];
endmodule

module inversebitpermute(input [63:0]a,output [63:0]b);
b[0]=a[63];b[1]=a[12];b[2]=a[25];b[3]=a[38];b[4]=a[51];b[5]=a[0];b[6]=a[13];b[7]=a[26];b[8]=a[39];b[9]=a[52];b[10]=a[1];b[11]=a[14];b[12]=a[27];b[13]=a[40];b[14]=a[53];b[15]=a[2];b[16]=a[15];b[17]=a[28];b[18]=a[41];b[19]=a[54];b[20]=a[3];b[21]=a[16];b[22]=a[29];b[23]=a[42];b[24]=a[55];b[25]=a[4];b[26]=a[17];b[27]=a[30];b[28]=a[43];b[29]=a[56];b[30]=a[5];b[31]=a[18];b[32]=a[31];b[33]=a[44];b[34]=a[57];b[35]=a[6];b[36]=a[19];b[37]=a[32];b[38]=a[45];b[39]=a[58];b[40]=a[7];b[41]=a[20];b[42]=a[33];b[43]=a[46];b[44]=a[59];b[45]=a[8];b[46]=a[21];b[47]=a[34];b[48]=a[47];b[49]=a[60];b[50]=a[9];b[51]=a[22];b[52]=a[35];b[53]=a[48];b[54]=a[61];b[55]=a[10];b[56]=a[23];b[57]=a[36];b[58]=a[49];b[59]=a[62];b[60]=a[11];b[61]=a[24];b[62]=a[37];b[63]=a[50];
endmodule
